module instruction_decode(	write_register, clock, reset,Reg2Loc, MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc,
						Branchreg, instruction, write_back, PC_branch_link_in, read_data1, read_data2,
						RegWrite_in, RegWrite_out, read_register1_out, read_register2_out, stall, PC_out_IF_ID, PC_mux, sign_extend_out,
						Uncondbranch);
input clock, reset, RegWrite_in, stall;
input [31:0] instruction;
input [4:0] write_register;
input [63:0] write_back, PC_branch_link_in, PC_out_IF_ID;

output [63:0] 	read_data1, read_data2, sign_extend_out, PC_mux;
output RegWrite_out, Reg2Loc, MemRead, MemtoReg, MemWrite, ALUSrc, 
				Uncondbranch, Branchreg;
output [1:0] ALUOp;
output [4:0] read_register1_out, read_register2_out;

//mux met Rd (instr[4:0]) en Rm (instr[20:16]) geschakeld door Reg2Loc
wire [4:0] read_register_2;
n_mux mux2(.in1(instruction[20:16]),.in2(instruction[4:0]),.out(read_register_2),.select(Reg2Loc));

//mux met write_back van MEM/WB pipeline register en PC_branch_link_in
//geschakeld door Branchlink
wire [63:0] write_data;
n_mux mux1(.in1(write_back),.in2(PC_branch_link_in),.out(write_data),.select(Branchlink));

assign read_register1_out = instruction[9:5];
assign read_register2_out = read_register_2;



//mux's voor stall
wire Reg2Loc_in, Branch_in, MemRead_in, MemtoReg_in, MemWrite_in, ALUSrc_in, RegWrite_in, Uncondbranch_in,
		Branchlink_in, Branchreg_in,Branchlink,Branch;				
n_mux n_mux_Reg2Loc(.in1(Reg2Loc_in), .in2(0), .out(Reg2Loc), .select(stall));
n_mux n_mux_Branch(.in1(Branch_in), .in2(0), .out(Branch), .select(stall));
n_mux n_mux_MemRead(.in1(MemRead_in), .in2(0), .out(MemRead), .select(stall));
n_mux n_mux_MemtoReg(.in1(MemtoReg_in), .in2(0), .out(MemtoReg), .select(stall));
n_mux n_mux_MemWrite(.in1(MemWrite_in), .in2(0), .out(MemWrite), .select(stall));
n_mux n_mux_ALUSrc(.in1(ALUSrc_in), .in2(0), .out(ALUSrc), .select(stall));
n_mux n_mux_RegWrite(.in1(RegWrite_in), .in2(0), .out(RegWrite_out), .select(stall));
n_mux n_mux_Uncondbranch(.in1(Uncondbranch_in), .in2(0), .out(Uncondbranch), .select(stall));
n_mux n_mux_Branchlink(.in1(Branchlink_in), .in2(0), .out(Branchlink), .select(stall));
n_mux n_mux_Branchreg(.in1(Branchreg_in), .in2(0), .out(Branchreg), .select(stall));

wire not_zero;
control control(.clock(clock), 
				.instruction(instruction[31:21]), 
				.Reg2Loc(Reg2Loc_in), 
				.Branch(Branch_in), 
				.MemRead(MemRead_in), 
				.MemtoReg(MemtoReg_in), 
				.ALUOp(ALUOp), 
				.MemWrite(MemWrite_in), 
				.ALUSrc(ALUSrc_in), 
				.RegWrite(RegWrite_in), 
				.Uncondbranch(Uncondbranch_in), 
				.Branchlink(Branchlink_in), 
				.Branchreg(Branchreg_in), 
				.not_zero(not_zero));
registers registers(.Read_register_1(instruction[9:5]), 
					.Read_register_2(read_register_2), 
					.Write_register(write_register), 
					.Write_data(write_data), 
					.RegWrite(RegWrite_in), 
					.Read_data_1(read_data1), 
					.Read_data_2(read_data2), 
					.clock(clock), 
					.reset(reset));
		
//bepaalde delen van de instructies sign extenden naar 64 bits
wire [63:0] sign_extend_out, shift_left_2_out, PC_CB, PC_mux, PC_mux_link;
sign_extend sign_extend(.in(instruction),.out(sign_extend_out));
shift_left_2 shift_left_2(sign_extend_out,shift_left_2_out);

//sign extended waarde offset optellen bij PC_out
alu_add add_pc_m(PC_out_IF_ID,shift_left_2_out,PC_CB);
			
wire alu_zero;					
n_mux mux_zero_not_zero(.in1(zero),.in2(!zero),.out(alu_zero),.select(not_zero));


wire or_out, and_out;
assign or_out = and_out | Uncondbranch;
assign and_out = Branch & alu_zero;
//selecteren tussen PC_inc en PC_CB
n_mux n_mux_PC_inc_CB(.in1(PC_out_IF_ID), .in2(PC_CB), .out(PC_mux), .select(or_out));

//kijken of read_data1 gelijk is aan 0
reg zero;
always @(read_data1) begin
	if (read_data1 == 64'b0) zero <= 1;
	else zero <= 0;
end

endmodule