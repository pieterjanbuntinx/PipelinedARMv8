module instruction_decode(	write_register, clock, reset,Reg2Loc, Branch, MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, Uncondbranch,
						Branchlink, Branchreg, not_zero, instruction, write_back, PC_branch_link_in, read_data1, read_data2, sign_extend_out,
						RegWrite_in, RegWrite_out, read_register1_out, read_register2_out, stall);
input clock, reset, RegWrite_in, stall;
input [31:0] instruction;
input [4:0] write_register;
input [63:0] write_back, PC_branch_link_in;

output [63:0] sign_extend_out, read_data1, read_data2,Reg2Loc, Branch, MemRead, MemtoReg, ALUOp, MemWrite, ALUSrc, Uncondbranch, Branchlink, Branchreg, not_zero;
output RegWrite_out;
output [4:0] read_register1_out, read_register2_out;

//mux met Rd (instr[4:0]) en Rm (instr[20:16]) geschakeld door Reg2Loc
wire [4:0] read_register_2;
n_mux mux2(.in1(instruction[20:16]),.in2(instruction[4:0]),.out(read_register_2),.select(Reg2Loc));

//mux met write_back van MEM/WB pipeline register en PC_branch_link_in
//geschakeld door Branchlink
wire [63:0] write_data;
n_mux mux1(.in1(write_back),.in2(PC_branch_link_in),.out(write_data),.select(Branchlink));

assign read_register1_out = instruction[9:5];
assign read_register2_out = read_register_2;

//mux's voor stall
wire Reg2Loc_in, Branch_in, MemRead_in, MemtoReg_in, MemWrite_in, ALUSrc_in, RegWrite_in, Uncondbranch_in,
		Branchlink_in, Branchreg_in;				
n_mux n_mux_Reg2Loc(.in1(Reg2Loc_in), .in2(0), .out(Reg2Loc), .select(stall));
n_mux n_mux_Branch(.in1(Branch_in), .in2(0), .out(Branch), .select(stall));
n_mux n_mux_MemRead(.in1(MemRead_in), .in2(0), .out(MemRead), .select(stall));
n_mux n_mux_MemtoReg(.in1(MemtoReg_in), .in2(0), .out(MemtoReg), .select(stall));
n_mux n_mux_MemWrite(.in1(MemWrite_in), .in2(0), .out(MemWrite), .select(stall));
n_mux n_mux_ALUSrc(.in1(ALUSrc_in), .in2(0), .out(ALUSrc), .select(stall));
n_mux n_mux_RegWrite(.in1(RegWrite_in), .in2(0), .out(RegWrite), .select(stall));
n_mux n_mux_Uncondbranch(.in1(Uncondbranch_in), .in2(0), .out(Uncondbranch), .select(stall));
n_mux n_mux_Branchlink(.in1(Branchlink_in), .in2(0), .out(Branchlink), .select(stall));
n_mux n_mux_Branchreg(.in1(Branchreg_in), .in2(0), .out(Branchreg), .select(stall));

control control(.clock(clock), 
				.instruction(instruction[31:21]), 
				.Reg2Loc(Reg2Loc_in), 
				.Branch(Branch_in), 
				.MemRead(MemRead_in), 
				.MemtoReg(MemtoReg_in), 
				.ALUOp(ALUOp), 
				.MemWrite(MemWrite_in), 
				.ALUSrc(ALUSrc_in), 
				.RegWrite(RegWrite_in), 
				.Uncondbranch(Uncondbranch_in), 
				.Branchlink(Branchlink_in), 
				.Branchreg(Branchreg_in), 
				.not_zero(not_zero));
registers registers(.Read_register_1(instruction[9:5]), 
					.Read_register_2(read_register_2), 
					.Write_register(write_register), 
					.Write_data(write_data), 
					.RegWrite(MEM_WB_RegWrite), 
					.Read_data_1(read_data1), 
					.Read_data_2(read_data2), 
					.clock(clock), 
					.reset(reset));

//bepaalde delen van de instructies sign extenden naar 64 bits
sign_extend sign_extend(.in(instruction),.out(sign_extend_out));

endmodule