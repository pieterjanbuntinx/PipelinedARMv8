module ID_EX(clock, reset, wren, PC_out_in, read_data1, read_data2, s_extended_in